/*
PBLM:Build a circuit with no inputs and one output that outputs a constant 0
*/
module constant_zero(
  output zero
);
  assign zero=1'b0;
endmodule
